`timescale 1ns / 1ps

module ALU_ctrl( funct, ALU_OP,ALU_CTRL );

    input [5:0] funct;
	input [1:0] ALU_OP;
    output [3:0]ALU_CTRL;
   
	
	
	
	   /* add your design */   
	


endmodule
